module tm1638(
    input clk,          // Входной тактовый сигнал
    input rst,          // Сигнал сброса

    input data_latch,   // Сигнал защелки для начала передачи данных
    inout [7:0] data,   // Двунаправленная шина данных
    input rw,           // Сигнал чтения/записи (1 - чтение, 0 - запись)

    output busy,        // Сигнал занятости модуля

    output sclk,        // Выходной тактовый сигнал для передачи данных
    input  dio_in,      // Входной сигнал данных
    output reg dio_out  // Выходной сигнал данных (добавлен reg)
    );

    // Локальные параметры для делителя тактовой частоты
    localparam CLK_DIV = 3;  // Делитель тактовой частоты (работает на 12 МГц с CLK_DIV = 3)
    localparam CLK_DIV1 = CLK_DIV - 1;

    // Состояния конечного автомата
    localparam [1:0]
        S_IDLE      = 2'h0,  // Состояние ожидания
        S_WAIT      = 2'h1,  // Состояние ожидания перед передачей
        S_TRANSFER  = 2'h2;  // Состояние передачи данных

    // Регистры для хранения текущего и следующего состояний
    reg [1:0] cur_state, next_state;

    // Регистры для управления тактовым сигналом
    reg [CLK_DIV1:0] sclk_d, sclk_q;

    // Регистры для хранения данных
    reg [7:0] data_d, data_q, data_out_d, data_out_q;

    // Регистры для управления выходным сигналом данных
    reg dio_out_d;

    // Счетчик для отслеживания переданных битов
    reg [2:0] ctr_d, ctr_q;

    // Управление двунаправленной шиной данных
    assign data = rw ? 8'hZZ : data_out_q;  // Если режим чтения, то шина в высокоимпедансном состоянии

    // Сигнал занятости: модуль занят, если не находится в состоянии ожидания
    assign busy = cur_state != S_IDLE;

    // Генерация тактового сигнала для передачи данных
    assign sclk = ~((~sclk_q[CLK_DIV1]) & (cur_state == S_TRANSFER));

    // Логика конечного автомата
    always @(*)
    begin
        // Инициализация значений по умолчанию
        sclk_d = sclk_q;
        data_d = data_q;
        dio_out_d = dio_out;
        ctr_d = ctr_q;
        data_out_d = data_out_q;
        next_state = cur_state;

        // Логика в зависимости от текущего состояния
        case(cur_state)
            S_IDLE: begin
                sclk_d = 0;  // Сброс тактового сигнала
                if (data_latch) begin  // Если активирована защелка
                    // Если режим чтения, сбросить данные, иначе зафиксировать данные для отправки
                    data_d = rw ? data : 8'b0;
                    next_state = S_WAIT;  // Переход в состояние ожидания
                end
            end

            S_WAIT: begin
                sclk_d = sclk_q + 4'd1;  // Увеличение счетчика тактового сигнала
                // Ожидание середины тактового импульса
                if (sclk_q == {1'b0, {CLK_DIV1{1'b1}}}) begin
                    sclk_d = 0;  // Сброс счетчика тактового сигнала
                    next_state = S_TRANSFER;  // Переход в состояние передачи данных
                end
            end

            S_TRANSFER: begin
                sclk_d = sclk_q + 4'd1;  // Увеличение счетчика тактового сигнала
                if (sclk_q == 0) begin
                    // Начало тактового импульса: вывод старшего бита данных
                    dio_out_d = data_q[0];

                end else if (sclk_q == {1'b0, {CLK_DIV1{1'b1}}}) begin
                    // Середина тактового импульса: чтение данных от устройства
                    data_d = {dio_in, data_q[7:1]};

                end else if (&sclk_q) begin
                    // Конец тактового импульса: увеличение счетчика битов
                    ctr_d = ctr_q + 3'd1;

                    if (&ctr_q) begin
                        // Если все биты переданы, переход в состояние ожидания
                        next_state = S_IDLE;
                        data_out_d = data_q;  // Сохранение полученных данных

                        dio_out_d = 0;  // Сброс выходного сигнала данных
                    end
                end
            end

            default:
                next_state = S_IDLE;  // По умолчанию переход в состояние ожидания
        endcase
    end

    // Блок обновления регистров на каждом такте
    always @(posedge clk)
    begin
        if (rst)  // Если активен сигнал сброса
        begin
            cur_state <= S_IDLE;  // Сброс состояния
            sclk_q <= 0;  // Сброс счетчика тактового сигнала
            ctr_q <= 0;  // Сброс счетчика битов
            dio_out <= 0;  // Сброс выходного сигнала данных
            data_q <= 0;  // Сброс регистра данных
            data_out_q <= 0;  // Сброс регистра выходных данных
        end
        else
        begin
            cur_state <= next_state;  // Обновление состояния
            sclk_q <= sclk_d;  // Обновление счетчика тактового сигнала
            ctr_q <= ctr_d;  // Обновление счетчика битов
            dio_out <= dio_out_d;  // Обновление выходного сигнала данных
            data_q <= data_d;  // Обновление регистра данных
            data_out_q <= data_out_d;  // Обновление регистра выходных данных
        end
    end
endmodule