module top(
    input clk,  // Входной тактовый сигнал

    output reg tm_cs,  // Выходной сигнал выбора чипа (Chip Select) для TM1638
    output tm_clk,     // Выходной тактовый сигнал для TM1638
    inout  tm_dio      // Двунаправленный сигнал данных для TM1638
    );

    // Локальные параметры для удобства чтения кода
    localparam 
        HIGH    = 1'b1,  // Логическая единица
        LOW     = 1'b0;  // Логический ноль

    // Локальные параметры для кодирования сегментов цифр на дисплее
    localparam [6:0]
        S_0     = 7'b0111111,  // Цифра 0                    3F
        S_1     = 7'b0000110,  // Цифра 1 7'b0000110         6
        S_2     = 7'b1011011,  // Цифра 2                    5B
        S_3     = 7'b1001111,  // Цифра 3                    4F
        S_4     = 7'b1100110,  // Цифра 4                    66
        S_5     = 7'b1101101,  // Цифра 5                    6D
        S_6     = 7'b1111101,  // Цифра 6                    7D
        S_7     = 7'b0000111,  // Цифра 7                    7
        S_8     = 7'b1111111,  // Цифра 8                    7F
        S_9     = 7'b1101111,  // Цифра 9                    6F
        S_BLK   = 7'b0000000;  // Пустой символ (все сегменты выключены)
/*
                       //hgfedcba             --a--
                      8'b00111111, // 0      |     |
                      8'b00000110, // 1      f     b      dcba
                      8'b01011011, // 2      |     |
                      8'b01001111, // 3       --g--
                      8'b01100110, // 4      |     |
                      8'b01101101, // 5      e     c
                      8'b01111101, // 6      |     |
                      8'b00000111};// 7       --d--
*/
    // Локальные параметры для команд управления TM1638
    localparam [7:0]
        C_READ  = 8'b01000010,  // Команда чтения данных  42
        C_WRITE = 8'b01000000,  // Команда записи данных  40
        C_DISP  = 8'b10001111,  // Команда включения дисплея с максимальной яркостью 8F
        C_ADDR  = 8'b11000000;  // Команда установки начального адреса   C0

    localparam CLK_DIV = 19;  // Скорость сканирования (делитель тактовой частоты)

    // Регистры для управления состоянием
    reg rst = HIGH;  // Регистр сброса
    reg [5:0] instruction_step;  // Текущий шаг выполнения инструкции
    reg [7:0] keys;  // Регистр для хранения состояния клавиш

    // Регистры для анимации "бегущего огня"
    reg [7:0] larson;  // Регистр для хранения состояния светодиодов
    reg larson_dir;    // Направление движения "бегущего огня"
    reg [CLK_DIV:0] counter;  // Счетчик для управления скоростью анимации

    // Настройка тристабильного вывода для дисплея
    //   tm_dio     - физический вывод
    //   dio_in     - для чтения данных с дисплея
    //   dio_out    - для отправки данных на дисплей
    //   tm_rw      - выбор режима (ввод/вывод)
    reg tm_rw;
    wire dio_in;  // Входной сигнал данных
    wire dio_out; // Выходной сигнал данных

    // Управление тристабильным выводом
    assign tm_dio = tm_rw ? dio_out : 1'bz;  // Если tm_rw = 1, то вывод данных, иначе высокоимпедансное состояние
    assign dio_in = tm_dio;  // Чтение данных с вывода

    /*
    SB_IO #(
        .PIN_TYPE(6'b101001),
        .PULLUP(1'b1)
    ) tm_dio_io (
        .PACKAGE_PIN(tm_dio),
        .OUTPUT_ENABLE(tm_rw),
        .D_IN_0(dio_in),
        .D_OUT_0(dio_out)
    );
    */

    // Настройка модуля TM1638 с тристабильным выводом
    //   tm_in      - данные, прочитанные с модуля
    //   tm_out     - данные, записываемые в модуль
    //   tm_latch   - сигнал защелки для чтения/записи данных
    //   tm_rw      - выбор режима (чтение/запись)
    //   busy       - сигнал занятости модуля
    //   tm_clk     - тактовый сигнал данных
    //   dio_in     - данные, прочитанные с дисплея
    //   dio_out    - данные, отправляемые на дисплей
    //   tm_data    - тристабильный вывод данных к модулю
    reg tm_latch;  // Сигнал защелки
    wire busy;     // Сигнал занятости модуля
    wire [7:0] tm_data, tm_in;  // Данные для обмена с модулем
    reg [7:0] tm_out;  // Данные для отправки на модуль

    assign tm_in = tm_data;  // Чтение данных с модуля
    assign tm_data = tm_rw ? tm_out : 8'hZZ;  // Управление тристабильным выводом

    // Подключение модуля TM1638
    tm1638 u_tm1638 (
        .clk(clk),
        .rst(rst),
        .data_latch(tm_latch),
        .data(tm_data),
        .rw(tm_rw),
        .busy(busy),
        .sclk(tm_clk),
        .dio_in(dio_in),
        .dio_out(dio_out)
    );

   

 // Задача для отображения цифры на дисплее
    task display_digit;
        input [2:0] key;  // Номер клавиши
        input [6:0] segs;  // Сегменты для отображения цифры

        begin
            tm_latch <= HIGH;  // Активировать защелку

            if (keys[key])
                tm_out <= {1'b1, S_BLK[6:0]};  // Включить десятичную точку
            else
                tm_out <= {1'b0, segs};  // Выключить десятичную точку
        end
    endtask



    // Задача для анимации светодиодов
    task display_led;
        input [2:0] dot;  // Номер светодиода

        begin
            tm_latch <= HIGH;  // Активировать защелку
            tm_out <= {7'b0, larson[dot]};  // Установить состояние светодиода
        end
    endtask

    // Основной блок, работающий на каждом положительном фронте тактового сигнала
    always @(posedge clk) begin
        if (rst) begin  // Если активен сигнал сброса
            instruction_step <= 6'b0;  // Сброс шага выполнения инструкции
            tm_cs <= HIGH;  // Деактивировать выбор чипа
            tm_rw <= HIGH;  // Установить режим записи
            rst <= LOW;  // Сбросить сигнал сброса

            counter <= 0;  // Сбросить счетчик
            keys <= 8'b0;  // Сбросить состояние клавиш
            larson_dir <= 0;  // Сбросить направление анимации
            larson <= 8'b00010000;  // Инициализировать состояние светодиодов

        end else begin
            if (&counter) begin  // Если счетчик достиг максимума
                larson_dir <= larson[6] ? 0 : larson[1] ? 1 : larson_dir;  // Изменить направление анимации

                if (larson_dir)
                    larson <= {larson[6:0], larson[7]};  // Сдвиг вправо
                else
                    larson <= {larson[0], larson[7:1]};  // Сдвиг влево
            end

            if (counter[0] && ~busy) begin  // Если счетчик кратен 2 и модуль не занят
                case (instruction_step)
                       // *** ЧТЕНИЕ КЛАВИШ ***
                    1:  {tm_cs, tm_rw}     <= {LOW, HIGH};  // Активировать выбор чипа и режим записи
                    2:  {tm_latch, tm_out} <= {HIGH, C_READ};  // Установить режим чтения
                    3:  {tm_latch, tm_rw}  <= {HIGH, LOW};  // Переключиться на режим чтения

                    // Чтение состояния клавиш S1 - S8
                    4:  {keys[7], keys[3]} <= {tm_in[0], tm_in[4]};  // Чтение первой пары клавиш
                    5:  {tm_latch}         <= {HIGH};  // Активировать защелку
                    6:  {keys[6], keys[2]} <= {tm_in[0], tm_in[4]};  // Чтение второй пары клавиш
                    7:  {tm_latch}         <= {HIGH};  // Активировать защелку
                    8:  {keys[5], keys[1]} <= {tm_in[0], tm_in[4]};  // Чтение третьей пары клавиш
                    9:  {tm_latch}         <= {HIGH};  // Активировать защелку
                    10: {keys[4], keys[0]} <= {tm_in[0], tm_in[4]};  // Чтение четвертой пары клавиш
                    11: {tm_cs}            <= {HIGH};  // Деактивировать выбор чипа

                    // *** ОТОБРАЖЕНИЕ НА ДИСПЛЕЕ ***
                    12: {tm_cs, tm_rw}     <= {LOW, HIGH};  // Активировать выбор чипа и режим записи
                    13: {tm_latch, tm_out} <= {HIGH, C_WRITE};  // Установить режим записи
                    14: {tm_cs}            <= {HIGH};  // Деактивировать выбор чипа

                    15: {tm_cs, tm_rw}     <= {LOW, HIGH};  // Активировать выбор чипа и режим записи
                    16: {tm_latch, tm_out} <= {HIGH, C_ADDR};  // Установить начальный адрес

                    17: display_digit(3'd7, S_1);  // Отобразить цифру 1
                    18: display_led(3'd0);        // Управление светодиодом 1

                    19: display_digit(3'd6, S_2);  // Отобразить цифру 2
                    20: display_led(3'd1);        // Управление светодиодом 2

                    21: display_digit(3'd5, S_3);  // Отобразить цифру 3
                    22: display_led(3'd2);        // Управление светодиодом 3

                    23: display_digit(3'd4, S_4);  // Отобразить цифру 4
                    24: display_led(3'd3);        // Управление светодиодом 4

                    25: display_digit(3'd3, S_5);  // Отобразить цифру 5
                    26: display_led(3'd4);        // Управление светодиодом 5

                    27: display_digit(3'd2, S_6);  // Отобразить цифру 6
                    28: display_led(3'd5);        // Управление светодиодом 6

                    29: display_digit(3'd1, S_7);  // Отобразить цифру 7
                    30: display_led(3'd6);        // Управление светодиодом 7

                    31: display_digit(3'd0, S_8);  // Отобразить цифру 8
                    32: display_led(3'd7);        // Управление светодиодом 8

                    33: {tm_cs}            <= {HIGH};  // Деактивировать выбор чипа

                    34: {tm_cs, tm_rw}     <= {LOW, HIGH};  // Активировать выбор чипа и режим записи
                    35: {tm_latch, tm_out} <= {HIGH, C_DISP};  // Включить дисплей с максимальной яркостью
                    36: {tm_cs, instruction_step} <= {HIGH, 6'b0};  // Деактивировать выбор чипа и сбросить шаг выполнения инструкции

                endcase

                instruction_step <= instruction_step + 6'd1;  // Переход к следующему шагу

            end else if (busy) begin  // Если модуль занят
                // Деактивировать защелку на следующем такте
                tm_latch <= LOW;
            end

            counter <= counter + 21'd1;  // Увеличение счетчика
        end
    end
endmodule